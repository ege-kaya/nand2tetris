`include "Mux16.v"

module Mux16_tb();

    reg [15:0] a;
    reg [15:0] b;
    reg sel;
    wire [15:0] out;

    initial begin

        $dumpfile("Mux16_tb.vcd");
        $dumpvars(0, Mux16_tb);

        a = 16'b0000000000000000; b = 16'b0000000000000000; sel = 0;
        #5 a = 16'b0000000000000000; b = 16'b1111111111111111; sel = 1;
        #5 a = 16'b0000000000000000; b = 16'b0001001000110100; sel = 0;
        #5 a = 16'b0000000000000000; b = 16'b0001001000110100; sel = 1;
        #5 a = 16'b1001100001110110; b = 16'b0000000000000000; sel = 0;
        #5 a = 16'b1001100001110110; b = 16'b0000000000000000; sel = 1;
        #5 a = 16'b1010101010101010; b = 16'b0101010101010101; sel = 0;
        #5 a = 16'b1010101010101010; b = 16'b0101010101010101; sel = 1;
        #5 $finish;

    end

    Mux16 U_Mux16(.out(out), .a(a), .b(b), .sel(sel));

endmodule
