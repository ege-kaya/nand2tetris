`include "Mux4Way16.v"

module Mux4Way16_tb();

    reg [15:0] a;
    reg [15:0] b;
    reg [15:0] c;
    reg [15:0] d;
    reg [1:0] sel;

    wire [15:0] out;

    initial begin

        $dumpfile("Mux4Way16_tb.vcd");
        $dumpvars(0, Mux4Way16_tb);

        a = 16'b0000000000000000; b = 16'b0000000000000000;
        c = 16'b0000000000000000; d = 16'b0000000000000000;
        sel = 2'b00;
        #5 a = 16'b0000000000000000; b = 16'b0000000000000000;
        c = 16'b0000000000000000; d = 16'b0000000000000000;
        sel = 2'b01;
        #5 a = 16'b0000000000000000; b = 16'b0000000000000000;
        c = 16'b0000000000000000; d = 16'b0000000000000000;
        sel = 2'b10;
        #5 a = 16'b0000000000000000; b = 16'b0000000000000000;
        c = 16'b0000000000000000; d = 16'b0000000000000000;
        sel = 2'b11;
        #5 a = 16'b0001001000110100; b = 16'b1001100001110110;
        c = 16'b1010101010101010; d = 16'b0101010101010101;
        sel = 2'b00;
        #5 a = 16'b0001001000110100; b = 16'b1001100001110110;
        c = 16'b1010101010101010; d = 16'b0101010101010101;
        sel = 2'b01;
        #5 a = 16'b0001001000110100; b = 16'b1001100001110110;
        c = 16'b1010101010101010; d = 16'b0101010101010101;
        sel = 2'b10;
        #5 a = 16'b0001001000110100; b = 16'b1001100001110110;
        c = 16'b1010101010101010; d = 16'b0101010101010101;
        sel = 2'b11;

        #5 $finish;

    end

    Mux4Way16 U_Mux4Way16(.out(out), .a(a), .b(b), .c(c), .d(d), .sel(sel));

endmodule
